module mux_4_1 (

input selo,

sell,

input 10,

il,

12,

13,

output wire y);

wire y0, yl;

mux_2_1 ml (sell, i2, 13, y1);

mux_2_1 m2 (sell, i0, il, y0);

mux_2_1 m3 (sel0, y0, y1, y);

endmodule

module mux_2_1 (

input sel,

input 10, il,

output y);

assign y = sel? il: 10;

endmodule
